module new();
endmodule
